`define _BUILD_TIME_H_ 32'h20250318
`define _BUILD_TIME_L_ 32'h092614
`define _SVN_VER_ 32'hUnversioned directory


