`define _BUILD_TIME_H_ 32'h20250207
`define _BUILD_TIME_L_ 32'h161808
`define _SVN_VER_ 32'hUnversioned directory

